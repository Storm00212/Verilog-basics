// This is a simple Verilog program that prints "Hello, World!" to the console.

module hello_world;

  initial begin
    $display("Hello, World!");
  end

endmodule
